
module test_beach(clk,rst);
input logic clk;
input logic rst;

simple_cpu simple_cpu_inst(clk,rst);
endmodule